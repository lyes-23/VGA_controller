library ieee; 
use ieee.std_logic_vector.all; 
use ieee.numeric_std.all;



entity affiche_obj is 
port(
x,y : in std_logic_vector(11 downto 0);